module pc_reg (
    ports
);
    
endmodule